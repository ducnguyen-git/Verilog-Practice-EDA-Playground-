module unsigned_mul_32bit_beha (HI, LO, A, B);
  // output list
  output [31:0] HI;
  output [31:0] LO;
  // input list
  input [31:0] A;
  input [31:0] B;
  
  reg [31:0] HI;
  reg [31:0] LO;
  
  always @(A or B) begin
    {HI,LO} = A * B;
  end  

endmodule